/**
 * PLL configuration
 *
 * This Verilog module was generated automatically
 * using the icepll tool from the IceStorm project.
 * Use at your own risk.
 *
 * Given input frequency:       100.000 MHz
 * Requested output frequency:   33.333 MHz
 * Achieved output frequency:    33.333 MHz
 */
`default_nettype none
module pll(
	input  wire in,
	output wire out,
	output wire reset
	);
	wire clk_out;
SB_PLL40_CORE #(
		.FEEDBACK_PATH("SIMPLE"),
		.DIVR(4'b1000),		// DIVR =  8
		.DIVF(7'b0101111),	// DIVF = 47
		.DIVQ(3'b100),		// DIVQ =  4
		.FILTER_RANGE(3'b001)	// FILTER_RANGE = 1
	) uut (
		.LOCK(reset),
		.RESETB(1'b1),
		.BYPASS(1'b0),
		.REFERENCECLK(in),
		.PLLOUTGLOBAL(clk_out)
		);
	
	SB_GB Clock_Buffer (
		.USER_SIGNAL_TO_GLOBAL_BUFFER (clk_out),
		.GLOBAL_BUFFER_OUTPUT (out)
	);

endmodule
